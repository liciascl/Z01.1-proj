library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity carrinho is
	port (
    x1, x2, x3, x4 : in  STD_LOGIC;
    y1, y2: out STD_LOGIC_VECTOR(1 downto 0));
end entity;

architecture arch of carrinho is

begin

end architecture;

-- Elementos de Sistemas
-- developed by Luciano Soares
-- file: CPU.vhd
-- date: 4/4/2017

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity CPU is
  port(
    clock:       in  STD_LOGIC;                        -- sinal de clock para CPU
    reset:       in  STD_LOGIC;                        -- reinicia toda a CPU (inclusive o Program Counter)
    inM:         in  STD_LOGIC_VECTOR(15 downto 0) := "0000000000000000";    -- dados lidos da memória RAM
    instruction: in  STD_LOGIC_VECTOR(17 downto 0) := "000000000000000000";    -- instrução (dados) vindos da memória ROM
    outM:        out STD_LOGIC_VECTOR(15 downto 0);    -- dados para gravar na memória RAM
    writeM:      out STD_LOGIC;                        -- faz a memória RAM gravar dados da entrada
    addressM:    out STD_LOGIC_VECTOR(14 downto 0);    -- envia endereço para a memória RAM
    pcout:       out STD_LOGIC_VECTOR(14 downto 0)     -- endereço para ser enviado a memória ROM
    );
end entity;

architecture arch of CPU is

  component Mux16 is
    port (
      a:   in  STD_LOGIC_VECTOR(15 downto 0);
      b:   in  STD_LOGIC_VECTOR(15 downto 0);
      sel: in  STD_LOGIC;
      q:   out STD_LOGIC_VECTOR(15 downto 0)
      );
  end component;

  component ALU is
    port (
      x,y:   in STD_LOGIC_VECTOR(15 downto 0);
      zx:    in STD_LOGIC;
      nx:    in STD_LOGIC;
      zy:    in STD_LOGIC;
      ny:    in STD_LOGIC;
      f:     in STD_LOGIC;
      no:    in STD_LOGIC;
      zr:    out STD_LOGIC;
      ng:    out STD_LOGIC;
      saida: out STD_LOGIC_VECTOR(15 downto 0)
      );
  end component;

  component Register16 is
    port(
      clock:   in std_logic;
      input:   in STD_LOGIC_VECTOR(15 downto 0);
      load:    in std_logic;
      output: out STD_LOGIC_VECTOR(15 downto 0)
      );
  end component;

  component pc is
    port(
      clock     : in  STD_LOGIC;
      increment : in  STD_LOGIC;
      load      : in  STD_LOGIC;
      reset     : in  STD_LOGIC;
      input     : in  STD_LOGIC_VECTOR(15 downto 0);
      output    : out STD_LOGIC_VECTOR(15 downto 0)
      );
  end component;

  signal c_muxALUI_A: STD_LOGIC := '0'; 
  signal c_muxAM: STD_LOGIC := '0'; 
  signal c_zx: STD_LOGIC := '0'; 
  signal c_nx: STD_LOGIC := '0';
  signal c_zy: STD_LOGIC := '0';
  signal c_ny: STD_LOGIC := '0';
  signal c_f: STD_LOGIC := '0';
  signal c_no: STD_LOGIC := '0';
  signal c_loadA: STD_LOGIC := '0';
  signal c_loadD: STD_LOGIC := '0';
  signal c_loadPC: STD_LOGIC := '0';
  signal c_zr: std_logic := '0'; 
  signal c_ng: std_logic := '0'; 

  signal s_muxALUI_Aout: STD_LOGIC_VECTOR(15 downto 0);
  signal s_muxAM_out: STD_LOGIC_VECTOR(15 downto 0);
  signal s_regAout: STD_LOGIC_VECTOR(15 downto 0);
  signal s_regDout: STD_LOGIC_VECTOR(15 downto 0);
  signal s_ALUout: STD_LOGIC_VECTOR(15 downto 0);

  signal s_pcout: STD_LOGIC_VECTOR(15 downto 0);

begin
  MuxALUI_A: Mux16 port map(s_ALUout,instruction(15 downto 0),c_muxALUI_A,s_muxALUI_Aout);  
  MuxAM: Mux16 port map(s_regAout,inM,c_muxAM,s_muxAM_out);  
  RegisterA: Register16 port map(clock,s_muxALUI_Aout,c_loadA,s_regAout);
  RegisterD: Register16 port map(clock,s_ALUout,c_loadD,s_regDout);
  ProgCont: pc port map(clock,'1',c_loadPC,reset,s_regAout,s_pcout);

  ula: ALU port map(s_regDout,s_muxAM_out,c_zx,c_nx,c_zy,c_ny,c_f,c_no,c_zr,c_ng,s_ALUout);
  outM <= s_ALUout;
  addressM <= s_regAout(14 downto 0);
  pcout <= s_pcout(14 downto 0);
  
  inst: process(instruction,c_ng,c_zr) is
  begin
  if instruction(17) = '0' then
  c_muxALUI_A <= '1';
  c_muxAM <= '0';
  c_zx <= '0';
  c_nx <= '0';
  c_zy <= '0';
  c_ny <= '0';
  c_f <= '0';
  c_no <= '0';
  c_loadA <= '1';
  c_loadD <= '0';
  writeM <= '0';
  c_loadPC <= '0';
  elsif instruction(17) = '1' then
  c_zx <= instruction(12);
  c_nx <= instruction(11);
  c_zy <= instruction(10);
  c_ny <= instruction(9);
  c_f <= instruction(8);
  c_no <= instruction(7);

  c_muxALUI_A <= '0';
  c_muxAM <= instruction(13);

  c_loadA <= instruction(3);
  c_loadD <= instruction(4);
  writeM <= instruction(5);
  
  if ((instruction(2 downto 0) = "111") or  
  (c_ng = '1' and instruction(2) = '1') or 
  (c_zr = '1' and instruction(1) = '1') or  
  (c_zr = '0' and c_ng = '0' and instruction(0) = '1') ) then
  c_loadPC <= '1';
  else
  c_loadPC <= '0';
  end if;
  end if;

  end process inst;

  
end;

